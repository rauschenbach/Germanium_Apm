Germanium amplifier
* SPICE2 - ��� ��������� ���������� ��� �������

* ����������
C1 2 IN 47u
C2 0 2 240p
C3 3 0 47u
C4 9 0 47u
C5 11 8 240p
C6 12 OUT 470u
C7 4 13 430p
D1 15 14 diod
Q1 5 2 6 MP41
Q2 4 8 6 mp41
Q3 11 5 4 GT404G
Q4 16 15 OUT GT404G
Q5 4 13 17 GT402G
Q6 4 17 18 GT806B
Q7 OUT 16 19 GT806B
R1 0 2 10k
R2 4 5 240
R3 3 6 8200
R4 7 3 8.2k
R5 9 8 1.2k
R6 8 OUT 33600
R7 11 13 51
R8 13 14 220.5
R9 12 15 1.8k
R10 7 12 1.8k
R11 OUT 17 15
R12 7 16 15
R13 OUT 18 1
R14 7 19 1
R15 0 OUT 8

* ���������
**V1 in 0 dc 0 ac 1 sin 0 0.5 5k
V1 in 0 dc 0 ac SIN 0 0.5 1K 0 0 

V2 7 0 dc 25 
V3 4 0 dc -25 

* ������
.MODEL MP41 PNP LEVEL=1 AF=1 BF=140 BR=4 CJC=90P CJE=30P CJS=0 EG=0.72 FC=500M
+ IKF=50M IKR=0 IRB=0.1M IS=3U ISC=0.6U ISE=.3U ITF=0 KF=0 MJC=0.5 MJE=0.5 MJS=0
+ NC=1.28 NE=1.28 NF=1 NR=1 PTF=0 RB=150 RBM=50 RC=0 RE=0 TF=0.1U TR=1.U VAF=15
+ VAR=0 VJC=750M VJE=750M VJS=750M VTF=0 XCJC=1 XTB=0 XTF=0 XTI=3

.MODEL GT404G NPN LEVEL=1 AF=1 BF=160 BR=9.4 CJC=2.86N CJE=2.08N CJS=0 EG=0.67
+ FC=500M IKF=2.5 IKR=200M IRB=0 IS=28U ISC=800N ISE=1.55U ITF=11.194M KF=0
+ MJC=3.5 MJE=4.05 MJS=0 NC=2 NE=2 NF=1.09 NR=1 PTF=0 RB=5 RBM=0 RC=100M RE=440M
+ TF=113N TR=448.17N VAF=35 VAR=0 VJC=750M VJE=750M VJS=750M VTF=10 XCJC=1 XTB=0
+ XTF=500M XTI=3

.MODEL diod D AF=1 BV=30 CJO=3.5PF EG=0.67 FC=500M IBV=1.00E-04 IS=8U KF=0
+ M=0.22 N=1.483 RS=1.85 TT=20N VJ=0.1 XTI=3

.MODEL GT402G PNP LEVEL=1 AF=1 BF=200 BR=9.5 CJC=580P CJE=400P CJS=0 EG=0.67
+ FC=500M IKF=3.5 IKR=500M IRB=0 IS=4.9U ISC=300N ISE=180N ITF=40.9U KF=0 MJC=3.9
+ MJE=5.7 MJS=0 NC=2 NE=1.9 NF=1.1 NR=1 PTF=0 RB=0 RBM=0 RC=200M RE=400M TF=75.56N
+ TR=96.58N VAF=18.3 VAR=0 VJC=850M VJE=850M VJS=750M VTF=10 XCJC=1 XTB=0 XTF=1.79
+ XTI=3

.MODEL GT806B PNP LEVEL=1 AF=1 BF=50 BR=1.000000004658M CJC=370.122683039208P
+ CJE=562.77720137022P CJS=0 EG=1.11 FC=500.000001073757M IKF=716.919946780524M
+ IKR=10.000001364568M IRB=0 IS=10.256643913003F ISC=98.557590750318P
+ ISE=.000000144458F ITF=63.387718169127F KF=0 MJC=383.692916282016M
+ MJE=483.990197021103M MJS=0 NC=2.000000003374 NE=650.541221795828M
+ NF=853.951123357701M NR=1 PTF=0 RB=0 RBM=0 RC=42.059429791057M
+ RE=92.22764856181M TF=20.342135167303N TR=999.999996592669M VAF=100 VAR=0
+ VJC=700.000000047339M VJE=750.097338903212M VJS=750M VTF=10.012794593207 XCJC=1
+ XTB=0 XTF=522.521126058016M XTI=3
*

.control
destroy all
tran 1u 5m .005m



setplot
setplot tran1 
plot  v(in) v(out) xlabel time[s]  ylabel 'In, Out [V]' 


ac dec 25 1Hz 100megHz 
setplot ac1 
set units = degrees
plot vp(out) 

let phase = unwrap(vp(out)) 
plot phase xlabel f[Hz] ylabel 'Magnitude[dB], Phase[deg]'


tran 100m 1 0 1
fourier 1 v(out)


.endc

.END


